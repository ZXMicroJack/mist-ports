module cos (
	x,
	y
);
	input [9:0] x;
	output wire [7:0] y;
	wire [2055:0] qcos = 2056'b111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111111011111110111111101111110011111100111111001111110011111100111111001111110011111100111110101111101011111010111110101111101011111010111110001111100011111000111110001111100011110110111101101111011011110110111101001111010011110100111101001111010011110010111100101111001011110010111100001111000011110000111011101110111011101110111011101110110011101100111011001110101011101010111010101110100011101000111010001110011011100110111001101110010011100100111001001110001011100010111000101110000011100000110111101101111011011110110111001101110011011010110110101101101011011000110110001101011011010110110101001101010011010100110100101101001011010000110100001100111011001110110011001100110011001010110010101100100011001000110001101100011011000100110001001100001011000010110000001100000010111110101111101011110010111100101110101011101010111000101110001011011010110110101101001011001010110010101100001011000010101110101011101010110010101010101010101010100010101000101001101010010010100100101000101010001010100000100111101001111010011100100111001001101010011000100110001001011010010100100101001001001010010000100100001000111010001110100011001000101010001010100010001000011010000110100001001000001010000010100000000111111001111100011111000111101001111000011110000111011001110100011101000111001001110000011100000110111001101100011010100110101001101000011001100110011001100100011000100110000001100000010111100101110001011010010110100101100001010110010101000101010001010010010100000100111001001110010011000100101001001000010010000100011001000100010000100100001001000000001111100011110000111100001110100011100000110110001101100011010000110010001100000011000000101110001011000010101000101000001010000010011000100100001000100010001000100000000111100001110000011010000110100001100000010110000101000001010000010010000100000000111000001100000011000000101000001000000001100000010000000100000000100000000;
	assign y = ((x >= 10'd0) && (x < 10'd257) ? 8'd128 + qcos[(256 - x) * 8+:8] : ((x >= 10'd257) && (x < 10'd513) ? 8'd128 - qcos[((256 - 10'd512) + x) * 8+:8] : ((x >= 10'd513) && (x < 10'd769) ? 8'd128 - qcos[((256 + 10'd512) - x) * 8+:8] : 8'd128 + qcos[(256 + x) * 8+:8])));
endmodule
