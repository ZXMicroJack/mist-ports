module lfsr(output wire[22:0] rnd);
   assign rnd = 23'haaa;
endmodule
